// Code your testbench here
// or browse Examples
module repeat_code;
  initial begin
    
    repeat(5)begin
      $display("this is repeat output ");
      $display("ur offerletter is coming soon");
      $display("------------------------------");
    end
  end
    endmodule
